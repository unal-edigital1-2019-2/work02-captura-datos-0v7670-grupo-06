`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:52:24 11/14/2019 
// Design Name: 
// Module Name:    captura_de_datos 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module captura_de_datos(VSYNC,HREF,HSYNC,a,
    );
output VSYNC,HREF,HSYNC,a;//declaracion
reg color [7:0];
endmodule
